// Control block for brief
module brief_ctrl (
  clk,
  rst,
  en,
  gaussian_done,
  patch,
  written,
  binary_string
);

// parameters
parameter BITS = 8;
parameter WIDTH = 7;
parameter PNUM = 256;
parameter PATCHLEN = 961*8;

// inputs
input clk;
input rst;
// a single bit signaling if calculation should be done, from fast
input en;
// recieve the done signal from gaussian, if done, start operating
input gaussian_done;
// recieve the patch
input [PATCHLEN-1:0] patch;


// outputs
// a signal showing calculation is done, can pass next point
output reg written;
// patchread addr
// final result
output reg [PNUM-1:0] binary_string;

// internal variables
wire [PNUM-1:0] comp_res;
//integer i = 0;
reg idx;
reg en_buf;

wire [BITS-1:0] p [0:30][0:30];
wire [BITS-1:0] x1 [0:PNUM-1];
wire [BITS-1:0] y1 [0:PNUM-1];
wire [BITS-1:0] x2 [0:PNUM-1];
wire [BITS-1:0] y2 [0:PNUM-1];

// Declare and initialize the pattern of the points (x1, y1, x2, y2)
wire [31:0] pos [0:256*4];
assign {pos[0], pos[1], pos[2], pos[3], pos[4], pos[5], pos[6], pos[7],
        pos[8], pos[9], pos[10], pos[11], pos[12], pos[13], pos[14], pos[15], 
        pos[16], pos[17], pos[18], pos[19], pos[20], pos[21], pos[22], pos[23], 
        pos[24], pos[25], pos[26], pos[27], pos[28], pos[29], pos[30], pos[31], 
        pos[32], pos[33], pos[34], pos[35], pos[36], pos[37], pos[38], pos[39], 
        pos[40], pos[41], pos[42], pos[43], pos[44], pos[45], pos[46], pos[47], 
        pos[48], pos[49], pos[50], pos[51], pos[52], pos[53], pos[54], pos[55], 
        pos[56], pos[57], pos[58], pos[59], pos[60], pos[61], pos[62], pos[63], 
        pos[64], pos[65], pos[66], pos[67], pos[68], pos[69], pos[70], pos[71], 
        pos[72], pos[73], pos[74], pos[75], pos[76], pos[77], pos[78], pos[79], 
        pos[80], pos[81], pos[82], pos[83], pos[84], pos[85], pos[86], pos[87], 
        pos[88], pos[89], pos[90], pos[91], pos[92], pos[93], pos[94], pos[95], 
        pos[96], pos[97], pos[98], pos[99], pos[100], pos[101], pos[102], pos[103], 
        pos[104], pos[105], pos[106], pos[107], pos[108], pos[109], pos[110], pos[111], 
        pos[112], pos[113], pos[114], pos[115], pos[116], pos[117], pos[118], pos[119], 
        pos[120], pos[121], pos[122], pos[123], pos[124], pos[125], pos[126], pos[127], 
        pos[128], pos[129], pos[130], pos[131], pos[132], pos[133], pos[134], pos[135], 
        pos[136], pos[137], pos[138], pos[139], pos[140], pos[141], pos[142], pos[143], 
        pos[144], pos[145], pos[146], pos[147], pos[148], pos[149], pos[150], pos[151], 
        pos[152], pos[153], pos[154], pos[155], pos[156], pos[157], pos[158], pos[159], 
        pos[160], pos[161], pos[162], pos[163], pos[164], pos[165], pos[166], pos[167], 
        pos[168], pos[169], pos[170], pos[171], pos[172], pos[173], pos[174], pos[175], 
        pos[176], pos[177], pos[178], pos[179], pos[180], pos[181], pos[182], pos[183], 
        pos[184], pos[185], pos[186], pos[187], pos[188], pos[189], pos[190], pos[191], 
        pos[192], pos[193], pos[194], pos[195], pos[196], pos[197], pos[198], pos[199], 
        pos[200], pos[201], pos[202], pos[203], pos[204], pos[205], pos[206], pos[207], 
        pos[208], pos[209], pos[210], pos[211], pos[212], pos[213], pos[214], pos[215], 
        pos[216], pos[217], pos[218], pos[219], pos[220], pos[221], pos[222], pos[223], 
        pos[224], pos[225], pos[226], pos[227], pos[228], pos[229], pos[230], pos[231], 
        pos[232], pos[233], pos[234], pos[235], pos[236], pos[237], pos[238], pos[239], 
        pos[240], pos[241], pos[242], pos[243], pos[244], pos[245], pos[246], pos[247], 
        pos[248], pos[249], pos[250], pos[251], pos[252], pos[253], pos[254], pos[255], 
        pos[256], pos[257], pos[258], pos[259], pos[260], pos[261], pos[262], pos[263], 
        pos[264], pos[265], pos[266], pos[267], pos[268], pos[269], pos[270], pos[271], 
        pos[272], pos[273], pos[274], pos[275], pos[276], pos[277], pos[278], pos[279], 
        pos[280], pos[281], pos[282], pos[283], pos[284], pos[285], pos[286], pos[287], 
        pos[288], pos[289], pos[290], pos[291], pos[292], pos[293], pos[294], pos[295], 
        pos[296], pos[297], pos[298], pos[299], pos[300], pos[301], pos[302], pos[303], 
        pos[304], pos[305], pos[306], pos[307], pos[308], pos[309], pos[310], pos[311], 
        pos[312], pos[313], pos[314], pos[315], pos[316], pos[317], pos[318], pos[319], 
        pos[320], pos[321], pos[322], pos[323], pos[324], pos[325], pos[326], pos[327], 
        pos[328], pos[329], pos[330], pos[331], pos[332], pos[333], pos[334], pos[335], 
        pos[336], pos[337], pos[338], pos[339], pos[340], pos[341], pos[342], pos[343], 
        pos[344], pos[345], pos[346], pos[347], pos[348], pos[349], pos[350], pos[351], 
        pos[352], pos[353], pos[354], pos[355], pos[356], pos[357], pos[358], pos[359], 
        pos[360], pos[361], pos[362], pos[363], pos[364], pos[365], pos[366], pos[367], 
        pos[368], pos[369], pos[370], pos[371], pos[372], pos[373], pos[374], pos[375], 
        pos[376], pos[377], pos[378], pos[379], pos[380], pos[381], pos[382], pos[383], 
        pos[384], pos[385], pos[386], pos[387], pos[388], pos[389], pos[390], pos[391], 
        pos[392], pos[393], pos[394], pos[395], pos[396], pos[397], pos[398], pos[399], 
        pos[400], pos[401], pos[402], pos[403], pos[404], pos[405], pos[406], pos[407], 
        pos[408], pos[409], pos[410], pos[411], pos[412], pos[413], pos[414], pos[415], 
        pos[416], pos[417], pos[418], pos[419], pos[420], pos[421], pos[422], pos[423], 
        pos[424], pos[425], pos[426], pos[427], pos[428], pos[429], pos[430], pos[431], 
        pos[432], pos[433], pos[434], pos[435], pos[436], pos[437], pos[438], pos[439], 
        pos[440], pos[441], pos[442], pos[443], pos[444], pos[445], pos[446], pos[447], 
        pos[448], pos[449], pos[450], pos[451], pos[452], pos[453], pos[454], pos[455], 
        pos[456], pos[457], pos[458], pos[459], pos[460], pos[461], pos[462], pos[463], 
        pos[464], pos[465], pos[466], pos[467], pos[468], pos[469], pos[470], pos[471], 
        pos[472], pos[473], pos[474], pos[475], pos[476], pos[477], pos[478], pos[479], 
        pos[480], pos[481], pos[482], pos[483], pos[484], pos[485], pos[486], pos[487], 
        pos[488], pos[489pos], pos[490], pos[491], pos[492], pos[493], pos[494], pos[495], 
        pos[496], pos[497], pos[498], pos[499], pos[500], pos[501], pos[502], pos[503], 
        pos[504], pos[505], pos[506], pos[507], pos[508], pos[509], pos[510], pos[511], 
        pos[512], pos[513], pos[514], pos[515], pos[516], pos[517], pos[518], pos[519], 
        pos[520], pos[521], pos[522], pos[523], pos[524], pos[525], pos[526], pos[527], 
        pos[528], pos[529], pos[530], pos[531], pos[532], pos[533], pos[534], pos[535], 
        pos[536], pos[537], pos[538], pos[539], pos[540], pos[541], pos[542], pos[543], 
        pos[544], pos[545], pos[546], pos[547], pos[548], pos[549], pos[550], pos[551], 
        pos[552], pos[553], pos[554], pos[555], pos[556], pos[557], pos[558], pos[559], 
        pos[560], pos[561], pos[562], pos[563], pos[564], pos[565], pos[566], pos[567], 
        pos[568], pos[569], pos[570], pos[571], pos[572], pos[573], pos[574], pos[575], 
        pos[576], pos[577], pos[578], pos[579], pos[580], pos[581], pos[582], pos[583], 
        pos[584], pos[585], pos[586], pos[587], pos[588], pos[589], pos[590], pos[591], 
        pos[592], pos[593], pos[594], pos[595], pos[596], pos[597], pos[598], pos[599], 
        pos[600], pos[601], pos[602], pos[603], pos[604], pos[605], pos[606], pos[607], 
        pos[608], pos[609], pos[610], pos[611], pos[612], pos[613], pos[614], pos[615], 
        pos[616], pos[617], pos[618], pos[619], pos[620], pos[621], pos[622], pos[623], 
        pos[624], pos[625], pos[626], pos[627], pos[628], pos[629], pos[630], pos[631], 
        pos[632], pos[633], pos[634], pos[635], pos[636], pos[637], pos[638], pos[639], 
        pos[640], pos[641], pos[642], pos[643], pos[644], pos[645], pos[646], pos[647], 
        pos[648], pos[649], pos[650], pos[651], pos[652], pos[653], pos[654], pos[655], 
        pos[656], pos[657], pos[658], pos[659], pos[660], pos[661], pos[662], pos[663], 
        pos[664], pos[665], pos[666], pos[667], pos[668], pos[669], pos[670], pos[671], 
        pos[672], pos[673], pos[674], pos[675], pos[676], pos[677], pos[678], pos[679], 
        pos[680], pos[681], pos[682], pos[683], pos[684], pos[685], pos[686], pos[687], 
        pos[688], pos[689], pos[690], pos[691], pos[692], pos[693], pos[694], pos[695], 
        pos[696], pos[697], pos[698], pos[699], pos[700], pos[701], pos[702], pos[703], 
        pos[704], pos[705], pos[706], pos[707], pos[708], pos[709], pos[710], pos[711], 
        pos[712], pos[713], pos[714], pos[715], pos[716], pos[717], pos[718], pos[719], 
        pos[720], pos[721], pos[722], pos[723], pos[724], pos[725], pos[726], pos[727], 
        pos[728], pos[729], pos[730], pos[731], pos[732], pos[733], pos[734], pos[735], 
        pos[736], pos[737], pos[738], pos[739], pos[740], pos[741], pos[742], pos[743], 
        pos[744], pos[745pos], pos[746], pos[747], pos[748], pos[749], pos[750], pos[751], 
        pos[752], pos[753], pos[754], pos[755], pos[756], pos[757], pos[758], pos[759], 
        pos[760], pos[761], pos[762], pos[763], pos[764], pos[765], pos[766], pos[767], 
        pos[768], pos[769], pos[770], pos[771], pos[772], pos[773], pos[774], pos[775], 
        pos[776], pos[777], pos[778], pos[779], pos[780], pos[781], pos[782], pos[783], 
        pos[784], pos[785], pos[786], pos[787], pos[788], pos[789], pos[790], pos[791], 
        pos[792], pos[793], pos[794], pos[795], pos[796], pos[797], pos[798], pos[799], 
        pos[800], pos[801], pos[802], pos[803], pos[804], pos[805], pos[806], pos[807], 
        pos[808], pos[809], pos[810], pos[811], pos[812], pos[813], pos[814], pos[815], 
        pos[816], pos[817], pos[818], pos[819], pos[820], pos[821], pos[822], pos[823], 
        pos[824], pos[825], pos[826], pos[827], pos[828], pos[829], pos[830], pos[831], 
        pos[832], pos[833], pos[834], pos[835], pos[836], pos[837], pos[838], pos[839], 
        pos[840], pos[841], pos[842], pos[843], pos[844], pos[845], pos[846], pos[847], 
        pos[848], pos[849], pos[850], pos[851], pos[852], pos[853], pos[854], pos[855], 
        pos[856], pos[857], pos[858], pos[859], pos[860], pos[861], pos[862], pos[863], 
        pos[864], pos[865], pos[866], pos[867], pos[868], pos[869], pos[870], pos[871], 
        pos[872], pos[873], pos[874], pos[875], pos[876], pos[877], pos[878], pos[879], 
        pos[880], pos[881], pos[882], pos[883], pos[884], pos[885], pos[886], pos[887], 
        pos[888], pos[889], pos[890], pos[891], pos[892], pos[893], pos[894], pos[895], 
        pos[896], pos[897], pos[898], pos[899], pos[900], pos[901], pos[902], pos[903], 
        pos[904], pos[905], pos[906], pos[907], pos[908], pos[909], pos[910], pos[911], 
        pos[912], pos[913], pos[914], pos[915], pos[916], pos[917], pos[918], pos[919], 
        pos[920], pos[921], pos[922], pos[923], pos[924], pos[925], pos[926], pos[927], 
        pos[928], pos[929], pos[930], pos[931], pos[932], pos[933], pos[934], pos[935], 
        pos[936], pos[937], pos[938], pos[939], pos[940], pos[941], pos[942], pos[943], 
        pos[944], pos[945], pos[946], pos[947], pos[948], pos[949], pos[950], pos[951], 
        pos[952], pos[953], pos[954], pos[955], pos[956], pos[957], pos[958], pos[959], 
        pos[960], pos[961], pos[962], pos[963], pos[964], pos[965], pos[966], pos[967], 
        pos[968], pos[969], pos[970], pos[971], pos[972], pos[973], pos[974], pos[975], 
        pos[976], pos[977], pos[978], pos[979], pos[980], pos[981], pos[982], pos[983], 
        pos[984], pos[985], pos[986], pos[987], pos[988], pos[989], pos[990], pos[991], 
        pos[992], pos[993], pos[994], pos[995], pos[996], pos[997], pos[998], pos[999], 
        pos[1000], pos[1001], pos[1002], pos[1003], pos[1004], pos[1005], pos[1006], pos[1007], 
        pos[1008], pos[1009], pos[1010], pos[1011], pos[1012], pos[1013], pos[1014], pos[1015], 
        pos[1016], pos[1017], pos[1018], pos[1019], pos[1020], pos[1021], pos[1022], pos[1023]}
         = {
                    32'd8, -32'd3, 32'd9, 32'd5/*mean (0), correlation (0)*/,
                    32'd4, 32'd2, 32'd7, -32'd12/*mean (1.12461e-05), correlation (0.0437584)*/,
                    -32'd11, 32'd9, -32'd8, 32'd2/*mean (3.37382e-05), correlation (0.0617409)*/,
                    32'd7, -32'd12, 32'd12, -32'd13/*mean (5.62303e-05), correlation (0.0636977)*/,
                    32'd2, -32'd13, 32'd2, 32'd12/*mean (0.000134953), correlation (0.085099)*/,
                    32'd1, -32'd7, 32'd1, 32'd6/*mean (0.000528565), correlation (0.0857175)*/,
                    -32'd2, -32'd10, -32'd2, -32'd4/*mean (0.0188821), correlation (0.0985774)*/,
                    -32'd13, -32'd13, -32'd11,-32'd8/*mean (0.0363135), correlation (0.0899616)*/,
                    -32'd13, -32'd3, -32'd12, -32'd9/*mean (0.121806), correlation (0.099849)*/,
                    32'd10, 32'd4, 32'd11, 32'd9/*mean (0.122065), correlation (0.093285)*/,
                    -32'd13, -32'd8, -32'd8, -32'd9/*mean (0.162787), correlation (0.0942748)*/,
                    -32'd11, 32'd7, -32'd9, 32'd12/*mean (0.21561), correlation (0.0974438)*/,
                    32'd7, 32'd7, 32'd12, 32'd6/*mean (0.160583), correlation (0.130064)*/,
                    -32'd4, -32'd5, -32'd3, 32'd0/*mean (0.228171), correlation (0.132998)*/,
                    -32'd13, 32'd2, -32'd12, -32'd3/*mean (0.00997526), correlation (0.145926)*/,
                    -32'd9, 32'd0, -32'd7, 32'd5/*mean (0.198234), correlation (0.143636)*/,
                    32'd12, -32'd6, 32'd12, -32'd1/*mean (0.0676226), correlation (0.16689)*/,
                    -32'd3, 32'd6, -32'd2, 32'd12/*mean (0.166847), correlation (0.171682)*/,
                    -32'd6, -32'd13, -32'd4,-32'd8/*mean (0.101215), correlation (0.179716)*/,
                    32'd11, -32'd13, 32'd12, -32'd8/*mean (0.200641), correlation (0.192279)*/,
                    32'd4, 32'd7, 32'd5, 32'd1/*mean (0.205106), correlation (0.186848)*/,
                    32'd5, -32'd3, 32'd10, -32'd3/*mean (0.234908), correlation (0.192319)*/,
                    32'd3, -32'd7, 32'd6, 32'd12/*mean (0.0709964), correlation (0.210872)*/,
                    -32'd8, -32'd7, -32'd6, -32'd2/*mean (0.0939834), correlation (0.212589)*/,
                    -32'd2, 32'd11, -32'd1, -32'd10/*mean (0.127778), correlation (0.20866)*/,
                    -32'd13, 32'd12, -32'd8, 32'd10/*mean (0.14783), correlation (0.206356)*/,
                    -32'd7, 32'd3, -32'd5, -32'd3/*mean (0.182141), correlation (0.198942)*/,
                    -32'd4, 32'd2, -32'd3, 32'd7/*mean (0.188237), correlation (0.21384)*/,
                    -32'd10, -32'd12, -32'd6, 32'd11/*mean (0.14865), correlation (0.23571)*/,
                    32'd5, -32'd12, 32'd6, -32'd7/*mean (0.222312), correlation (0.23324)*/,
                    32'd5, -32'd6, 32'd7,-32'd1/*mean (0.229082), correlation (0.23389)*/,
                    32'd1, 32'd0, 32'd4, -32'd5/*mean (0.241577), correlation (0.215286)*/,
                    32'd9, 32'd11, 32'd11, -32'd13/*mean (0.00338507), correlation (0.251373)*/,
                    32'd4, 32'd7, 32'd4, 32'd12/*mean (0.131005), correlation (0.257622)*/,
                    32'd2, -32'd1, 32'd4, 32'd4/*mean (0.152755), correlation (0.255205)*/,
                    -32'd4, -32'd12, -32'd2, 32'd7/*mean (0.182771), correlation (0.244867)*/,
                    -32'd8, -32'd5, -32'd7, -32'd10/*mean (0.186898), correlation (0.23901)*/,
                    32'd4, 32'd11, 32'd9, 32'd12/*mean (0.226226), correlation (0.258255)*/,
                    32'd0, -32'd8, 32'd1, -32'd13/*mean (0.0897886), correlation (0.274827)*/,
                    -32'd13, -32'd2, -32'd8, 32'd2/*mean (0.148774), correlation (0.28065)*/,
                    -32'd3, -32'd2, -32'd2, 32'd3/*mean (0.153048), correlation (0.283063)*/,
                    -32'd6, 32'd9, -32'd4, -32'd9/*mean (0.169523), correlation (0.278248)*/,
                    32'd8, 32'd12, 32'd10, 32'd7/*mean (0.225337), correlation (0.282851)*/,
                    32'd0, 32'd9, 32'd1, 32'd3/*mean (0.226687), correlation (0.278734)*/,
                    32'd7, -32'd5, 32'd11, -32'd10/*mean (0.00693882), correlation (0.305161)*/,
                    -32'd13, -32'd6, -32'd11, 32'd0/*mean (0.0227283), correlation (0.300181)*/,
                    32'd10, 32'd7, 32'd12, 32'd1/*mean (0.125517), correlation (0.31089)*/,
                    -32'd6, -32'd3, -32'd6, 32'd12/*mean (0.131748), correlation (0.312779)*/,
                    32'd10, -32'd9, 32'd12, -32'd4/*mean (0.144827), correlation (0.292797)*/,
                    -32'd13, 32'd8, -32'd8, -32'd12/*mean (0.149202), correlation (0.308918)*/,
                    -32'd13, 32'd0, -32'd8, -32'd4/*mean (0.160909), correlation (0.310013)*/,
                    32'd3, 32'd3, 32'd7, 32'd8/*mean (0.177755), correlation (0.309394)*/,
                    32'd5, 32'd7, 32'd10, -32'd7/*mean (0.212337), correlation (0.310315)*/,
                    -32'd1, 32'd7, 32'd1, -32'd12/*mean (0.214429), correlation (0.311933)*/,
                    32'd3, -32'd10, 32'd5, 32'd6/*mean (0.235807), correlation (0.313104)*/,
                    32'd2, -32'd4, 32'd3, -32'd10/*mean (0.00494827), correlation (0.344948)*/,
                    -32'd13, 32'd0, -32'd13, 32'd5/*mean (0.0549145), correlation (0.344675)*/,
                    -32'd13, -32'd7, -32'd12, 32'd12/*mean (0.103385), correlation (0.342715)*/,
                    -32'd13, 32'd3, -32'd11, 32'd8/*mean (0.134222), correlation (0.322922)*/,
                    -32'd7, 32'd12, -32'd4, 32'd7/*mean (0.153284), correlation (0.337061)*/,
                    32'd6, -32'd10, 32'd12, 32'd8/*mean (0.154881), correlation (0.329257)*/,
                    -32'd9, -32'd1, -32'd7, -32'd6/*mean (0.200967), correlation (0.33312)*/,
                    -32'd2, -32'd5, 32'd0, 32'd12/*mean (0.201518), correlation (0.340635)*/,
                    -32'd12, 32'd5, -32'd7, 32'd5/*mean (0.207805), correlation (0.335631)*/,
                    32'd3, -32'd10, 32'd8, -32'd13/*mean (0.224438), correlation (0.34504)*/,
                    -32'd7, -32'd7, -32'd4, 32'd5/*mean (0.239361), correlation (0.338053)*/,
                    -32'd3, -32'd2, -32'd1, -32'd7/*mean (0.240744), correlation (0.344322)*/,
                    32'd2, 32'd9, 32'd5, -32'd11/*mean (0.242949), correlation (0.34145)*/,
                    -32'd11, -32'd13, -32'd5, -32'd13/*mean (0.244028), correlation (0.336861)*/,
                    -32'd1, 32'd6, 32'd0,-32'd1/*mean (0.247571), correlation (0.343684)*/,
                    32'd5, -32'd3, 32'd5, 32'd2/*mean (0.000697256), correlation (0.357265)*/,
                    -32'd4, -32'd13, -32'd4, 32'd12/*mean (0.00213675), correlation (0.373827)*/,
                    -32'd9, -32'd6, -32'd9, 32'd6/*mean (0.0126856), correlation (0.373938)*/,
                    -32'd12, -32'd10, -32'd8, -32'd4/*mean (0.0152497), correlation (0.364237)*/,
                    32'd10, 32'd2, 32'd12, -32'd3/*mean (0.0299933), correlation (0.345292)*/,
                    32'd7, 32'd12, 32'd12, 32'd12/*mean (0.0307242), correlation (0.366299)*/,
                    -32'd7, -32'd13, -32'd6, 32'd5/*mean (0.0534975), correlation (0.368357)*/,
                    -32'd4, 32'd9, -32'd3, 32'd4/*mean (0.099865), correlation (0.372276)*/,
                    32'd7, -32'd1, 32'd12, 32'd2/*mean (0.117083), correlation (0.364529)*/,
                    -32'd7, 32'd6, -32'd5, 32'd1/*mean (0.126125), correlation (0.369606)*/,
                    -32'd13, 32'd11, -32'd12, 32'd5/*mean (0.130364), correlation (0.358502)*/,
                    -32'd3, 32'd7, -32'd2,-32'd6/*mean (0.131691), correlation (0.375531)*/,
                    32'd7, -32'd8, 32'd12, -32'd7/*mean (0.160166), correlation (0.379508)*/,
                    -32'd13, -32'd7, -32'd11, -32'd12/*mean (0.167848), correlation (0.353343)*/,
                    32'd1, -32'd3, 32'd12, 32'd12/*mean (0.183378), correlation (0.371916)*/,
                    32'd2, -32'd6, 32'd3, 32'd0/*mean (0.228711), correlation (0.371761)*/,
                    -32'd4, 32'd3, -32'd2, -32'd13/*mean (0.247211), correlation (0.364063)*/,
                    -32'd1, -32'd13, 32'd1, 32'd9/*mean (0.249325), correlation (0.378139)*/,
                    32'd7, 32'd1, 32'd8,-32'd6/*mean (0.000652272), correlation (0.411682)*/,
                    32'd1, -32'd1, 32'd3, 32'd12/*mean (0.00248538), correlation (0.392988)*/,
                    32'd9, 32'd1, 32'd12, 32'd6/*mean (0.0206815), correlation (0.386106)*/,
                    -32'd1, -32'd9, -32'd1, 32'd3/*mean (0.0364485), correlation (0.410752)*/,
                    -32'd13, -32'd13, -32'd10, 32'd5/*mean (0.0376068), correlation (0.398374)*/,
                    32'd7, 32'd7, 32'd10, 32'd12/*mean (0.0424202), correlation (0.405663)*/,
                    32'd12, -32'd5, 32'd12, 32'd9/*mean (0.0942645), correlation (0.410422)*/,
                    32'd6, 32'd3, 32'd7, 32'd11/*mean (0.1074), correlation (0.413224)*/,
                    32'd5, -32'd13, 32'd6, 32'd10/*mean (0.109256), correlation (0.408646)*/,
                    32'd2, -32'd12, 32'd2, 32'd3/*mean (0.131691), correlation (0.416076)*/,
                    32'd3, 32'd8, 32'd4, -32'd6/*mean (0.165081), correlation (0.417569)*/,
                    32'd2, 32'd6, 32'd12, -32'd13/*mean (0.171874), correlation (0.408471)*/,
                    32'd9, -32'd12, 32'd10, 32'd3/*mean (0.175146), correlation (0.41296)*/,
                    -32'd8, 32'd4, -32'd7, 32'd9/*mean (0.183682), correlation (0.402956)*/,
                    -32'd11, 32'd12, -32'd4, -32'd6/*mean (0.184672), correlation (0.416125)*/,
                    32'd1, 32'd12, 32'd2, -32'd8/*mean (0.191487), correlation (0.386696)*/,
                    32'd6, -32'd9, 32'd7, -32'd4/*mean (0.192668), correlation (0.394771)*/,
                    32'd2, 32'd3, 32'd3, -32'd2/*mean (0.200157), correlation (0.408303)*/,
                    32'd6, 32'd3, 32'd11, 32'd0/*mean (0.204588), correlation (0.411762)*/,
                    32'd3, -32'd3, 32'd8, -32'd8/*mean (0.205904), correlation (0.416294)*/,
                    32'd7, 32'd8, 32'd9, 32'd3/*mean (0.213237), correlation (0.409306)*/,
                    -32'd11, -32'd5, -32'd6, -32'd4/*mean (0.243444), correlation (0.395069)*/,
                    -32'd10, 32'd11, -32'd5, 32'd10/*mean (0.247672), correlation (0.413392)*/,
                    -32'd5, -32'd8, -32'd3, 32'd12/*mean (0.24774), correlation (0.411416)*/,
                    -32'd10, 32'd5, -32'd9, 32'd0/*mean (0.00213675), correlation (0.454003)*/,
                    32'd8, -32'd1, 32'd12, -32'd6/*mean (0.0293635), correlation (0.455368)*/,
                    32'd4, -32'd6, 32'd6, -32'd11/*mean (0.0404971), correlation (0.457393)*/,
                    -32'd10, 32'd12, -32'd8, 32'd7/*mean (0.0481107), correlation (0.448364)*/,
                    32'd4, -32'd2, 32'd6, 32'd7/*mean (0.050641), correlation (0.455019)*/,
                    -32'd2, 32'd0, -32'd2, 32'd12/*mean (0.0525978), correlation (0.44338)*/,
                    -32'd5, -32'd8, -32'd5, 32'd2/*mean (0.0629667), correlation (0.457096)*/,
                    32'd7, -32'd6, 32'd10, 32'd12/*mean (0.0653846), correlation (0.445623)*/,
                    -32'd9, -32'd13, -32'd8, -32'd8/*mean (0.0858749), correlation (0.449789)*/,
                    -32'd5, -32'd13, -32'd5, -32'd2/*mean (0.122402), correlation (0.450201)*/,
                    32'd8, -32'd8, 32'd9, -32'd13/*mean (0.125416), correlation (0.453224)*/,
                    -32'd9, -32'd11, -32'd9, 32'd0/*mean (0.130128), correlation (0.458724)*/,
                    32'd1, -32'd8, 32'd1, -32'd2/*mean (0.132467), correlation (0.440133)*/,
                    32'd7, -32'd4, 32'd9, 32'd1/*mean (0.132692), correlation (0.454)*/,
                    -32'd2, 32'd1, -32'd1, -32'd4/*mean (0.135695), correlation (0.455739)*/,
                    32'd11, -32'd6, 32'd12, -32'd11/*mean (0.142904), correlation (0.446114)*/,
                    -32'd12, -32'd9, -32'd6, 32'd4/*mean (0.146165), correlation (0.451473)*/,
                    32'd3, 32'd7, 32'd7, 32'd12/*mean (0.147627), correlation (0.456643)*/,
                    32'd5, 32'd5, 32'd10, 32'd8/*mean (0.152901), correlation (0.455036)*/,
                    32'd0, -32'd4, 32'd2, 32'd8/*mean (0.167083), correlation (0.459315)*/,
                    -32'd9, 32'd12, -32'd5, -32'd13/*mean (0.173234), correlation (0.454706)*/,
                    32'd0, 32'd7, 32'd2, 32'd12/*mean (0.18312), correlation (0.433855)*/,
                    -32'd1, 32'd2, 32'd1, 32'd7/*mean (0.185504), correlation (0.443838)*/,
                    32'd5, 32'd11, 32'd7, -32'd9/*mean (0.185706), correlation (0.451123)*/,
                    32'd3, 32'd5, 32'd6, -32'd8/*mean (0.188968), correlation (0.455808)*/,
                    -32'd13, -32'd4, -32'd8, 32'd9/*mean (0.191667), correlation (0.459128)*/,
                    -32'd5, 32'd9, -32'd3, -32'd3/*mean (0.193196), correlation (0.458364)*/,
                    -32'd4, -32'd7, -32'd3, -32'd12/*mean (0.196536), correlation (0.455782)*/,
                    32'd6, 32'd5, 32'd8, 32'd0/*mean (0.1972), correlation (0.450481)*/,
                    -32'd7, 32'd6, -32'd6, 32'd12/*mean (0.199438), correlation (0.458156)*/,
                    -32'd13, 32'd6, -32'd5, -32'd2/*mean (0.211224), correlation (0.449548)*/,
                    32'd1, -32'd10, 32'd3, 32'd10/*mean (0.211718), correlation (0.440606)*/,
                    32'd4, 32'd1, 32'd8, -32'd4/*mean (0.213034), correlation (0.443177)*/,
                    -32'd2, -32'd2, 32'd2, -32'd13/*mean (0.234334), correlation (0.455304)*/,
                    32'd2, -32'd12, 32'd12, 32'd12/*mean (0.235684), correlation (0.443436)*/,
                    -32'd2, -32'd13, 32'd0, -32'd6/*mean (0.237674), correlation (0.452525)*/,
                    32'd4, 32'd1, 32'd9, 32'd3/*mean (0.23962), correlation (0.444824)*/,
                    -32'd6, -32'd10, -32'd3, -32'd5/*mean (0.248459), correlation (0.439621)*/,
                    -32'd3, -32'd13, -32'd1, 32'd1/*mean (0.249505), correlation (0.456666)*/,
                    32'd7, 32'd5, 32'd12, -32'd11/*mean (0.00119208), correlation (0.495466)*/,
                    32'd4, -32'd2, 32'd5, -32'd7/*mean (0.00372245), correlation (0.484214)*/,
                    -32'd13, 32'd9, -32'd9, -32'd5/*mean (0.00741116), correlation (0.499854)*/,
                    32'd7, 32'd1, 32'd8, 32'd6/*mean (0.0208952), correlation (0.499773)*/,
                    32'd7, -32'd8, 32'd7, 32'd6/*mean (0.0220085), correlation (0.501609)*/,
                    -32'd7, -32'd4, -32'd7, 32'd1/*mean (0.0233806), correlation (0.496568)*/,
                    -32'd8, 32'd11, -32'd7, -32'd8/*mean (0.0236505), correlation (0.489719)*/,
                    -32'd13, 32'd6, -32'd12, -32'd8/*mean (0.0268781), correlation (0.503487)*/,
                    32'd2, 32'd4, 32'd3, 32'd9/*mean (0.0323324), correlation (0.501938)*/,
                    32'd10, -32'd5, 32'd12, 32'd3/*mean (0.0399235), correlation (0.494029)*/,
                    -32'd6, -32'd5, -32'd6, 32'd7/*mean (0.0420153), correlation (0.486579)*/,
                    32'd8, -32'd3, 32'd9, -32'd8/*mean (0.0548021), correlation (0.484237)*/,
                    32'd2, -32'd12, 32'd2, 32'd8/*mean (0.0616622), correlation (0.496642)*/,
                    -32'd11, -32'd2, -32'd10, 32'd3/*mean (0.0627755), correlation (0.498563)*/,
                    -32'd12, -32'd13, -32'd7, -32'd9/*mean (0.0829622), correlation (0.495491)*/,
                    -32'd11, 32'd0, -32'd10, -32'd5/*mean (0.0843342), correlation (0.487146)*/,
                    32'd5, -32'd3, 32'd11, 32'd8/*mean (0.0929937), correlation (0.502315)*/,
                    -32'd2, -32'd13, -32'd1, 32'd12/*mean (0.113327), correlation (0.48941)*/,
                    -32'd1, -32'd8, 32'd0, 32'd9/*mean (0.132119), correlation (0.467268)*/,
                    -32'd13, -32'd11, -32'd12, -32'd5/*mean (0.136269), correlation (0.498771)*/,
                    -32'd10, -32'd2, -32'd10, 32'd11/*mean (0.142173), correlation (0.498714)*/,
                    -32'd3, 32'd9, -32'd2,-32'd13/*mean (0.144141), correlation (0.491973)*/,
                    32'd2, -32'd3, 32'd3, 32'd2/*mean (0.14892), correlation (0.500782)*/,
                    -32'd9, -32'd13, -32'd4, 32'd0/*mean (0.150371), correlation (0.498211)*/,
                    -32'd4, 32'd6, -32'd3, -32'd10/*mean (0.152159), correlation (0.495547)*/,
                    -32'd4, 32'd12, -32'd2,-32'd7/*mean (0.156152), correlation (0.496925)*/,
                    -32'd6, -32'd11, -32'd4, 32'd9/*mean (0.15749), correlation (0.499222)*/,
                    32'd6, -32'd3, 32'd6, 32'd11/*mean (0.159211), correlation (0.503821)*/,
                    -32'd13, 32'd11, -32'd5, 32'd5/*mean (0.162427), correlation (0.501907)*/,
                    32'd11, 32'd11, 32'd12, 32'd6/*mean (0.16652), correlation (0.497632)*/,
                    32'd7, -32'd5, 32'd12, -32'd2/*mean (0.169141), correlation (0.484474)*/,
                    -32'd1, 32'd12, 32'd0, 32'd7/*mean (0.169456), correlation (0.495339)*/,
                    -32'd4, -32'd8, -32'd3, -32'd2/*mean (0.171457), correlation (0.487251)*/,
                    -32'd7, 32'd1, -32'd6, 32'd7/*mean (0.175), correlation (0.500024)*/,
                    -32'd13, -32'd12, -32'd8, -32'd13/*mean (0.175866), correlation (0.497523)*/,
                    -32'd7, -32'd2, -32'd6, -32'd8/*mean (0.178273), correlation (0.501854)*/,
                    -32'd8, 32'd5, -32'd6, -32'd9/*mean (0.181107), correlation (0.494888)*/,
                    -32'd5, -32'd1, -32'd4, 32'd5/*mean (0.190227), correlation (0.482557)*/,
                    -32'd13, 32'd7, -32'd8, 32'd10/*mean (0.196739), correlation (0.496503)*/,
                    32'd1, 32'd5, 32'd5, -32'd13/*mean (0.19973), correlation (0.499759)*/,
                    32'd1, 32'd0, 32'd10, -32'd13/*mean (0.204465), correlation (0.49873)*/,
                    32'd9, 32'd12, 32'd10, -32'd1/*mean (0.209334), correlation (0.49063)*/,
                    32'd5, -32'd8, 32'd10, -32'd9/*mean (0.211134), correlation (0.503011)*/,
                    -32'd1, 32'd11, 32'd1, -32'd13/*mean (0.212), correlation (0.499414)*/,
                    -32'd9, -32'd3, -32'd6, 32'd2/*mean (0.212168), correlation (0.480739)*/,
                    -32'd1, -32'd10, 32'd1, 32'd12/*mean (0.212731), correlation (0.502523)*/,
                    -32'd13, 32'd1, -32'd8, -32'd10/*mean (0.21327), correlation (0.489786)*/,
                    32'd8, -32'd11, 32'd10, -32'd6/*mean (0.214159), correlation (0.488246)*/,
                    32'd2, -32'd13, 32'd3, -32'd6/*mean (0.216993), correlation (0.50287)*/,
                    32'd7, -32'd13, 32'd12, -32'd9/*mean (0.223639), correlation (0.470502)*/,
                    -32'd10, -32'd10, -32'd5, -32'd7/*mean (0.224089), correlation (0.500852)*/,
                    -32'd10, -32'd8, -32'd8, -32'd13/*mean (0.228666), correlation (0.502629)*/,
                    32'd4, -32'd6, 32'd8, 32'd5/*mean (0.22906), correlation (0.498305)*/,
                    32'd3, 32'd12, 32'd8, -32'd13/*mean (0.233378), correlation (0.503825)*/,
                    -32'd4, 32'd2, -32'd3, -32'd3/*mean (0.234323), correlation (0.476692)*/,
                    32'd5, -32'd13, 32'd10, -32'd12/*mean (0.236392), correlation (0.475462)*/,
                    32'd4, -32'd13, 32'd5, -32'd1/*mean (0.236842), correlation (0.504132)*/,
                    -32'd9, 32'd9, -32'd4, 32'd3/*mean (0.236977), correlation (0.497739)*/,
                    32'd0, 32'd3, 32'd3, -32'd9/*mean (0.24314), correlation (0.499398)*/,
                    -32'd12, 32'd1, -32'd6, 32'd1/*mean (0.243297), correlation (0.489447)*/,
                    32'd3, 32'd2, 32'd4, -32'd8/*mean (0.00155196), correlation (0.553496)*/,
                    -32'd10, -32'd10, -32'd10, 32'd9/*mean (0.00239541), correlation (0.54297)*/,
                    32'd8, -32'd13, 32'd12, 32'd12/*mean (0.0034413), correlation (0.544361)*/,
                    -32'd8, -32'd12, -32'd6, -32'd5/*mean (0.003565), correlation (0.551225)*/,
                    32'd2, 32'd2, 32'd3, 32'd7/*mean (0.00835583), correlation (0.55285)*/,
                    32'd10, 32'd6, 32'd11, -32'd8/*mean (0.00885065), correlation (0.540913)*/,
                    32'd6, 32'd8, 32'd8, -32'd12/*mean (0.0101552), correlation (0.551085)*/,
                    -32'd7, 32'd10, -32'd6, 32'd5/*mean (0.0102227), correlation (0.533635)*/,
                    -32'd3, -32'd9, -32'd3, 32'd9/*mean (0.0110211), correlation (0.543121)*/,
                    -32'd1, -32'd13, -32'd1, 32'd5/*mean (0.0113473), correlation (0.550173)*/,
                    -32'd3, -32'd7, -32'd3, 32'd4/*mean (0.0140913), correlation (0.554774)*/,
                    -32'd8, -32'd2, -32'd8, 32'd3/*mean (0.017049), correlation (0.55461)*/,
                    32'd4, 32'd2, 32'd12, 32'd12/*mean (0.01778), correlation (0.546921)*/,
                    32'd2, -32'd5, 32'd3, 32'd11/*mean (0.0224022), correlation (0.549667)*/,
                    32'd6, -32'd9, 32'd11, -32'd13/*mean (0.029161), correlation (0.546295)*/,
                    32'd3, -32'd1, 32'd7, 32'd12/*mean (0.0303081), correlation (0.548599)*/,
                    32'd11, -32'd1, 32'd12, 32'd4/*mean (0.0355151), correlation (0.523943)*/,
                    -32'd3, 32'd0, -32'd3, 32'd6/*mean (0.0417904), correlation (0.543395)*/,
                    32'd4, -32'd11, 32'd4, 32'd12/*mean (0.0487292), correlation (0.542818)*/,
                    32'd2, -32'd4, 32'd2, 32'd1/*mean (0.0575124), correlation (0.554888)*/,
                    -32'd10, -32'd6, -32'd8, 32'd1/*mean (0.0594242), correlation (0.544026)*/,
                    -32'd13, 32'd7, -32'd11, 32'd1/*mean (0.0597391), correlation (0.550524)*/,
                    -32'd13, 32'd12, -32'd11, -32'd13/*mean (0.0608974), correlation (0.55383)*/,
                    32'd6, 32'd0, 32'd11, -32'd13/*mean (0.065126), correlation (0.552006)*/,
                    32'd0, -32'd1, 32'd1, 32'd4/*mean (0.074224), correlation (0.546372)*/,
                    -32'd13, 32'd3, -32'd9, -32'd2/*mean (0.0808592), correlation (0.554875)*/,
                    -32'd9, 32'd8, -32'd6, -32'd3/*mean (0.0883378), correlation (0.551178)*/,
                    -32'd13, -32'd6, -32'd8, -32'd2/*mean (0.0901035), correlation (0.548446)*/,
                    32'd5, -32'd9, 32'd8, 32'd10/*mean (0.0949843), correlation (0.554694)*/,
                    32'd2, 32'd7, 32'd3, -32'd9/*mean (0.0994152), correlation (0.550979)*/,
                    -32'd1, -32'd6, -32'd1, -32'd1/*mean (0.10045), correlation (0.552714)*/,
                    32'd9, 32'd5, 32'd11, -32'd2/*mean (0.100686), correlation (0.552594)*/,
                    32'd11, -32'd3, 32'd12, -32'd8/*mean (0.101091), correlation (0.532394)*/,
                    32'd3, 32'd0, 32'd3, 32'd5/*mean (0.101147), correlation (0.525576)*/,pos
                    -32'd1, 32'd4, 32'd0, 32'd10/*mean (0.105263), correlation (0.531498)*/,
                    32'd3, -32'd6, 32'd4, 32'd5/*mean (0.110785), correlation (0.540491)*/,
                    -32'd13, 32'd0, -32'd10, 32'd5/*mean (0.112798), correlation (0.536582)*/,
                    32'd5, 32'd8, 32'd12, 32'd11/*mean (0.114181), correlation (0.555793)*/,
                    32'd8, 32'd9, 32'd9, -32'd6/*mean (0.117431), correlation (0.553763)*/,
                    32'd7, -32'd4, 32'd8, -32'd12/*mean (0.118522), correlation (0.553452)*/,
                    -32'd10, 32'd4, -32'd10, 32'd9/*mean (0.12094), correlation (0.554785)*/,
                    32'd7, 32'd3, 32'd12, 32'd4/*mean (0.122582), correlation (0.555825)*/,
                    32'd9, -32'd7, 32'd10, -32'd2/*mean (0.124978), correlation (0.549846)*/,
                    32'd7, 32'd0, 32'd12, -32'd2/*mean (0.127002), correlation (0.537452)*/,
                    -32'd1, -32'd6, 32'd0, -32'd11/*mean (0.127148), correlation (0.547401)*/
            };


assign {p[0][0],  p[0][1],  p[0][2],  p[0][3],  p[0][4],  p[0][5],  p[0][6],  p[0][7], 
        p[0][8],  p[0][9],  p[0][10], p[0][11], p[0][12], p[0][13], p[0][14], p[0][15], 
        p[0][16], p[0][17], p[0][18], p[0][19], p[0][20], p[0][21], p[0][22], p[0][23], 
        p[0][24], p[0][25], p[0][26], p[0][27], p[0][28], p[0][29], p[0][30],
        p[1][0],  p[1][1],  p[1][2],  p[1][3],  p[1][4],  p[1][5],  p[1][6],  p[1][7], 
        p[1][8],  p[1][9],  p[1][10], p[1][11], p[1][12], p[1][13], p[1][14], p[1][15], 
        p[1][16], p[1][17], p[1][18], p[1][19], p[1][20], p[1][21], p[1][22], p[1][23], 
        p[1][24], p[1][25], p[1][26], p[1][27], p[1][28], p[1][29], p[1][30],
        p[2][0],  p[2][1],  p[2][2],  p[2][3],  p[2][4],  p[2][5],  p[2][6],  p[2][7], 
        p[2][8],  p[2][9],  p[2][10], p[2][11], p[2][12], p[2][13], p[2][14], p[2][15], 
        p[2][16], p[2][17], p[2][18], p[2][19], p[2][20], p[2][21], p[2][22], p[2][23], 
        p[2][24], p[2][25], p[2][26], p[2][27], p[2][28], p[2][29], p[2][30],
        p[3][0],  p[3][1],  p[3][2],  p[3][3],  p[3][4],  p[3][5],  p[3][6],  p[3][7], 
        p[3][8],  p[3][9],  p[3][10], p[3][11], p[3][12], p[3][13], p[3][14], p[3][15], 
        p[3][16], p[3][17], p[3][18], p[3][19], p[3][20], p[3][21], p[3][22], p[3][23], 
        p[3][24], p[3][25], p[3][26], p[3][27], p[3][28], p[3][29], p[3][30],
        p[4][0],  p[4][1],  p[4][2],  p[4][3],  p[4][4],  p[4][5],  p[4][6],  p[4][7], 
        p[4][8],  p[4][9],  p[4][10], p[4][11], p[4][12], p[4][13], p[4][14], p[4][15], 
        p[4][16], p[4][17], p[4][18], p[4][19], p[4][20], p[4][21], p[4][22], p[4][23], 
        p[4][24], p[4][25], p[4][26], p[4][27], p[4][28], p[4][29], p[4][30],
        p[5][0],  p[5][1],  p[5][2],  p[5][3],  p[5][4],  p[5][5],  p[5][6],  p[5][7], 
        p[5][8],  p[5][9],  p[5][10], p[5][11], p[5][12], p[5][13], p[5][14], p[5][15], 
        p[5][16], p[5][17], p[5][18], p[5][19], p[5][20], p[5][21], p[5][22], p[5][23], 
        p[5][24], p[5][25], p[5][26], p[5][27], p[5][28], p[5][29], p[5][30],
        p[6][0],  p[6][1],  p[6][2],  p[6][3],  p[6][4],  p[6][5],  p[6][6],  p[6][7], 
        p[6][8],  p[6][9],  p[6][10], p[6][11], p[6][12], p[6][13], p[6][14], p[6][15], 
        p[6][16], p[6][17], p[6][18], p[6][19], p[6][20], p[6][21], p[6][22], p[6][23], 
        p[6][24], p[6][25], p[6][26], p[6][27], p[6][28], p[6][29], p[6][30],
        p[7][0],  p[7][1],  p[7][2],  p[7][3],  p[7][4],  p[7][5],  p[7][6],  p[7][7], 
        p[7][8],  p[7][9],  p[7][10], p[7][11], p[7][12], p[7][13], p[7][14], p[7][15], 
        p[7][16], p[7][17], p[7][18], p[7][19], p[7][20], p[7][21], p[7][22], p[7][23], 
        p[7][24], p[7][25], p[7][26], p[7][27], p[7][28], p[7][29], p[7][30],
        p[8][0],  p[8][1],  p[8][2],  p[8][3],  p[8][4],  p[8][5],  p[8][6],  p[8][7], 
        p[8][8],  p[8][9],  p[8][10], p[8][11], p[8][12], p[8][13], p[8][14], p[8][15], 
        p[8][16], p[8][17], p[8][18], p[8][19], p[8][20], p[8][21], p[8][22], p[8][23], 
        p[8][24], p[8][25], p[8][26], p[8][27], p[8][28], p[8][29], p[8][30],
        p[9][0],  p[9][1],  p[9][2],  p[9][3],  p[9][4],  p[9][5],  p[9][6],  p[9][7], 
        p[9][8],  p[9][9],  p[9][10], p[9][11], p[9][12], p[9][13], p[9][14], p[9][15], 
        p[9][16], p[9][17], p[9][18], p[9][19], p[9][20], p[9][21], p[9][22], p[9][23], 
        p[9][24], p[9][25], p[9][26], p[9][27], p[9][28], p[9][29], p[9][30],
        p[10][0],  p[10][1],  p[10][2],  p[10][3],  p[10][4],  p[10][5],  p[10][6],  p[10][7], 
        p[10][8],  p[10][9],  p[10][10], p[10][11], p[10][12], p[10][13], p[10][14], p[10][15], 
        p[10][16], p[10][17], p[10][18], p[10][19], p[10][20], p[10][21], p[10][22], p[10][23], 
        p[10][24], p[10][25], p[10][26], p[10][27], p[10][28], p[10][29], p[10][30],
        p[11][0],  p[11][1],  p[11][2],  p[11][3],  p[11][4],  p[11][5],  p[11][6],  p[11][7], 
        p[11][8],  p[11][9],  p[11][10], p[11][11], p[11][12], p[11][13], p[11][14], p[11][15], 
        p[11][16], p[11][17], p[11][18], p[11][19], p[11][20], p[11][21], p[11][22], p[11][23], 
        p[11][24], p[11][25], p[11][26], p[11][27], p[11][28], p[11][29], p[11][30],
        p[12][0],  p[12][1],  p[12][2],  p[12][3],  p[12][4],  p[12][5],  p[12][6],  p[12][7], 
        p[12][8],  p[12][9],  p[12][10], p[12][11], p[12][12], p[12][13], p[12][14], p[12][15], 
        p[12][16], p[12][17], p[12][18], p[12][19], p[12][20], p[12][21], p[12][22], p[12][23], 
        p[12][24], p[12][25], p[12][26], p[12][27], p[12][28], p[12][29], p[12][30],
        p[13][0],  p[13][1],  p[13][2],  p[13][3],  p[13][4],  p[13][5],  p[13][6],  p[13][7], 
        p[13][8],  p[13][9],  p[13][10], p[13][11], p[13][12], p[13][13], p[13][14], p[13][15], 
        p[13][16], p[13][17], p[13][18], p[13][19], p[13][20], p[13][21], p[13][22], p[13][23], 
        p[13][24], p[13][25], p[13][26], p[13][27], p[13][28], p[13][29], p[13][30],
        p[14][0],  p[14][1],  p[14][2],  p[14][3],  p[14][4],  p[14][5],  p[14][6],  p[14][7], pos
        p[14][8],  p[14][9],  p[14][10], p[14][11], p[14][12], p[14][13], p[14][14], p[14][15], 
        p[14][16], p[14][17], p[14][18], p[14][19], p[14][20], p[14][21], p[14][22], p[14][23], 
        p[14][24], p[14][25], p[14][26], p[14][27], p[14][28], p[14][29], p[14][30],
        p[15][0],  p[15][1],  p[15][2],  p[15][3],  p[15][4],  p[15][5],  p[15][6],  p[15][7], 
        p[15][8],  p[15][9],  p[15][10], p[15][11], p[15][12], p[15][13], p[15][14], p[15][15], 
        p[15][16], p[15][17], p[15][18], p[15][19], p[15][20], p[15][21], p[15][22], p[15][23], 
        p[15][24], p[15][25], p[15][26], p[15][27], p[15][28], p[15][29], p[15][30],
        p[16][0],  p[16][1],  p[16][2],  p[16][3],  p[16][4],  p[16][5],  p[16][6],  p[16][7], 
        p[16][8],  p[16][9],  p[16][10], p[16][11], p[16][12], p[16][13], p[16][14], p[16][15], 
        p[16][16], p[16][17], p[16][18], p[16][19], p[16][20], p[16][21], p[16][22], p[16][23], 
        p[16][24], p[16][25], p[16][26], p[16][27], p[16][28], p[16][29], p[16][30],
        p[17][0],  p[17][1],  p[17][2],  p[17][3],  p[17][4],  p[17][5],  p[17][6],  p[17][7], 
        p[17][8],  p[17][9],  p[17][10], p[17][11], p[17][12], p[17][13], p[17][14], p[17][15], 
        p[17][16], p[17][17], p[17][18], p[17][19], p[17][20], p[17][21], p[17][22], p[17][23], 
        p[17][24], p[17][25], p[17][26], p[17][27], p[17][28], p[17][29], p[17][30],
        p[18][0],  p[18][1],  p[18][2],  p[18][3],  p[18][4],  p[18][5],  p[18][6],  p[18][7], 
        p[18][8],  p[18][9],  p[18][10], p[18][11], p[18][12], p[18][13], p[18][14], p[18][15], 
        p[18][16], p[18][17], p[18][18], p[18][19], p[18][20], p[18][21], p[18][22], p[18][23], 
        p[18][24], p[18][25], p[18][26], p[18][27], p[18][28], p[18][29], p[18][30],
        p[19][0],  p[19][1],  p[19][2],  p[19][3],  p[19][4],  p[19][5],  p[19][6],  p[19][7], 
        p[19][8],  p[19][9],  p[19][10], p[19][11], p[19][12], p[19][13], p[19][14], p[19][15], 
        p[19][16], p[19][17], p[19][18], p[19][19], p[19][20], p[19][21], p[19][22], p[19][23], 
        p[19][24], p[19][25], p[19][26], p[19][27], p[19][28], p[19][29], p[19][30],
        p[20][0],  p[20][1],  p[20][2],  p[20][3],  p[20][4],  p[20][5],  p[20][6],  p[20][7], 
        p[20][8],  p[20][9],  p[20][10], p[20][11], p[20][12], p[20][13], p[20][14], p[20][15], 
        p[20][16], p[20][17], p[20][18], p[20][19], p[20][20], p[20][21], p[20][22], p[20][23], 
        p[20][24], p[20][25], p[20][26], p[20][27], p[20][28], p[20][29], p[20][30],
        p[21][0],  p[21][1],  p[21][2],  p[21][3],  p[21][4],  p[21][5],  p[21][6],  p[21][7], 
        p[21][8],  p[21][9],  p[21][10], p[21][11], p[21][12], p[21][13], p[21][14], p[21][15], 
        p[21][16], p[21][17], p[21][18], p[21][19], p[21][20], p[21][21], p[21][22], p[21][23], 
        p[21][24], p[21][25], p[21][26], p[21][27], p[21][28], p[21][29], p[21][30],
        p[22][0],  p[22][1],  p[22][2],  p[22][3],  p[22][4],  p[22][5],  p[22][6],  p[22][7], 
        p[22][8],  p[22][9],  p[22][10], p[22][11], p[22][12], p[22][13], p[22][14], p[22][15], 
        p[22][16], p[22][17], p[22][18], p[22][19], p[22][20], p[22][21], p[22][22], p[22][23], 
        p[22][24], p[22][25], p[22][26], p[22][27], p[22][28], p[22][29], p[22][30],
        p[23][0],  p[23][1],  p[23][2],  p[23][3],  p[23][4],  p[23][5],  p[23][6],  p[23][7], 
        p[23][8],  p[23][9],  p[23][10], p[23][11], p[23][12], p[23][13], p[23][14], p[23][15], 
        p[23][16], p[23][17], p[23][18], p[23][19], p[23][20], p[23][21], p[23][22], p[23][23], 
        p[23][24], p[23][25], p[23][26], p[23][27], p[23][28], p[23][29], p[23][30],
        p[24][0],  p[24][1],  p[24][2],  p[24][3],  p[24][4],  p[24][5],  p[24][6],  p[24][7], 
        p[24][8],  p[24][9],  p[24][10], p[24][11], p[24][12], p[24][13], p[24][14], p[24][15], 
        p[24][16], p[24][17], p[24][18], p[24][19], p[24][20], p[24][21], p[24][22], p[24][23], 
        p[24][24], p[24][25], p[24][26], p[24][27], p[24][28], p[24][29], p[24][30],
        p[25][0],  p[25][1],  p[25][2],  p[25][3],  p[25][4],  p[25][5],  p[25][6],  p[25][7], 
        p[25][8],  p[25][9],  p[25][10], p[25][11], p[25][12], p[25][13], p[25][14], p[25][15], 
        p[25][16], p[25][17], p[25][18], p[25][19], p[25][20], p[25][21], p[25][22], p[25][23], 
        p[25][24], p[25][25], p[25][26], p[25][27], p[25][28], p[25][29], p[25][30],
        p[26][0],  p[26][1],  p[26][2],  p[26][3],  p[26][4],  p[26][5],  p[26][6],  p[26][7], 
        p[26][8],  p[26][9],  p[26][10], p[26][11], p[26][12], p[26][13], p[26][14], p[26][15], 
        p[26][16], p[26][17], p[26][18], p[26][19], p[26][20], p[26][21], p[26][22], p[26][23], 
        p[26][24], p[26][25], p[26][26], p[26][27], p[26][28], p[26][29], p[26][30],
        p[27][0],  p[27][1],  p[27][2],  p[27][3],  p[27][4],  p[27][5],  p[27][6],  p[27][7], 
        p[27][8],  p[27][9],  p[27][10], p[27][11], p[27][12], p[27][13], p[27][14], p[27][15], 
        p[27][16], p[27][17], p[27][18], p[27][19], p[27][20], p[27][21], p[27][22], p[27][23], 
        p[27][24], p[27][25], p[27][26], p[27][27], p[27][28], p[27][29], p[27][30],
        p[28][0],  p[28][1],  p[28][2],  p[28][3],  p[28][4],  p[28][5],  p[28][6],  p[28][7], 
        p[28][8],  p[28][9],  p[28][10], p[28][11], p[28][12], p[28][13], p[28][14], p[28][15], 
        p[28][16], p[28][17], p[28][18], p[28][19], p[28][20], p[28][21], p[28][22], p[28][23], 
        p[28][24], p[28][25], p[28][26], p[28][27], p[28][28], p[28][29], p[28][30],
        p[29][0],  p[29][1],  p[29][2],  p[29][3],  p[29][4],  p[29][5],  p[29][6],  p[29][7], 
        p[29][8],  p[29][9],  p[29][10], p[29][11], p[29][12], p[29][13], p[29][14], p[29][15], 
        p[29][16], p[29][17], p[29][18], p[29][19], p[29][20], p[29][21], p[29][22], p[29][23], 
        p[29][24], p[29][25], p[29][26], p[29][27], p[29][28], p[29][29], p[29][30],
        p[30][0],  p[30][1],  p[30][2],  p[30][3],  p[30][4],  p[30][5],  p[30][6],  p[30][7], 
        p[30][8],  p[30][9],  p[30][10], p[30][11], p[30][12], p[30][13], p[30][14], p[30][15], 
        p[30][16], p[30][17], p[30][18], p[30][19], p[30][20], p[30][21], p[30][22], p[30][23], 
        p[30][24], p[30][25], p[30][26], p[30][27], p[30][28], p[30][29], p[30][30]
        } = patch;

// generate 256 binary comparisons
genvar j;
generate
  for (j = 0; j<PNUM; j=j+1) begin
    assign x1[j] = pos[4*j]+15;
    assign y1[j] = pos[4*j+1]+15;
    assign x2[j] = pos[4*j+2]+15;
    assign y2[j] = pos[4*j+3]+15;
  end
endgenerate


genvar i;
generate
  for (i = 0; i<PNUM; i=i+1) begin
    binary_test bt (.x(p[y1[i]][x1[i]]),
                    .y(p[y2[i]][x2[i]]),
                    .result(comp_res[i]));
    /*binary_test bt (.x(patch[8*(481-pos[4*i]+31*pos[4*i+1]):8*(481-pos[4*i]+31*pos[4*i+1])-7]),
                    .y(patch[8*(481-pos[4*i+2]+31*pos[4*i+3]):8*(481-pos[4*i+2]+31*pos[4*i+3])-7]),
                    .result(comp_res[i]));*/
                    
  end
endgenerate



always @(posedge clk) begin
  en_buf <= en;
  if ((!rst) & en_buf & gaussian_done) begin
    binary_string <= comp_res;
    written <= 1'b1;
  end
  else begin
    binary_string <= 255'b0;
    written <= 1'b0;
  end 
end

  
endmodule
