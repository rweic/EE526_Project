module gaussian (
  // inputs
  input [391:0] input_pixels,
  // outputs
  output [7:0] result
);

// internal variables
reg [7:0] A [0:6][0:6];
integer i,j;
//integer result = 0;

// 7 * 7 mask
real mask [0:6][0:6];
/*mask = 
  {0.0049,    0.0092,    0.0134,    0.0152,    0.0134,    0.0092,    0.0049,
   0.0092,    0.0172,    0.0250,    0.0283,    0.0250,    0.0172,    0.0092,
   0.0134,    0.0250,    0.0364,    0.0412,    0.0364,    0.0250,    0.0134,
   0.0152,    0.0283,    0.0412,    0.0467,    0.0412,    0.0283,    0.0152,
   0.0134,    0.0250,    0.0364,    0.0412,    0.0364,    0.0250,    0.0134,
   0.0092,    0.0172,    0.0250,    0.0283,    0.0250,    0.0172,    0.0092,
   0.0049,    0.0092,    0.0134,    0.0152,    0.0134,    0.0092,    0.0049};*/

always@(input_pixels)
  begin
    {A[0][0],A[0][1],A[0][2],A[0][3],A[0][4],A[0][5],A[0][6],
     A[1][0],A[1][1],A[1][2],A[1][3],A[1][4],A[1][5],A[1][6],
     A[2][0],A[2][1],A[2][2],A[2][3],A[2][4],A[2][5],A[2][6],
     A[3][0],A[3][1],A[3][2],A[3][3],A[3][4],A[3][5],A[3][6],
     A[4][0],A[4][1],A[4][2],A[4][3],A[4][4],A[4][5],A[4][6],
     A[5][0],A[5][1],A[5][2],A[5][3],A[5][4],A[5][5],A[5][6],
     A[6][0],A[6][1],A[6][2],A[6][3],A[6][4],A[6][5],A[6][6]} <= input_pixels;
     
     
  end

endmodule
