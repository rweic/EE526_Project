module gaussian_core (
  clk,
  input_pixels,
  result
);

// parameters
parameter BITS = 8;
parameter WIDTH = 7;

// inputs
input clk;
input [391:0] input_pixels;
// outputs
output reg [7:0] result;

// Declare the gaussian mask
// wire [BITS-1:0] M[0:WIDTH-1][0:WIDTH-1];
wire [BITS-1:0] M [0:3][0:3];
assign {M[0][0],M[0][1],M[0][2],M[0][3],
        M[1][0],M[1][1],M[1][2],M[1][3],
        M[2][0],M[2][1],M[2][2],M[2][3],
        M[3][0],M[3][1],M[3][2],M[3][3]}
          = {8'd5,  8'd9,  8'd14, 8'd16,
             8'd9,  8'd18, 8'd26, 8'd29,
             8'd14, 8'd26, 8'd37, 8'd42,
             8'd16, 8'd29, 8'd42, 8'd28};

// internal variables
// reg [BITS-1:0] A [0:WIDTH-1][0:WIDTH-1];
wire [BITS-1:0] A [0:WIDTH-1][0:WIDTH-1];
//integer i,j;
//integer sum;
        
assign {A[0][0],A[0][1],A[0][2],A[0][3],A[0][4],A[0][5],A[0][6],
        A[1][0],A[1][1],A[1][2],A[1][3],A[1][4],A[1][5],A[1][6],
        A[2][0],A[2][1],A[2][2],A[2][3],A[2][4],A[2][5],A[2][6],
        A[3][0],A[3][1],A[3][2],A[3][3],A[3][4],A[3][5],A[3][6],
        A[4][0],A[4][1],A[4][2],A[4][3],A[4][4],A[4][5],A[4][6],
        A[5][0],A[5][1],A[5][2],A[5][3],A[5][4],A[5][5],A[5][6],
        A[6][0],A[6][1],A[6][2],A[6][3],A[6][4],A[6][5],A[6][6]} = input_pixels;

reg [17:0] prod [0:3][0:3];
always@(*) begin
  prod[0][0] <= M[0][0] * (A[0][0] + A[6][0] + A[0][6] + A[6][6]);
  prod[0][1] <= M[0][1] * (A[0][1] + A[6][1] + A[0][5] + A[6][5]);
  prod[0][2] <= M[0][2] * (A[0][2] + A[6][2] + A[0][4] + A[6][4]);
  prod[1][0] <= M[1][0] * (A[1][0] + A[5][0] + A[1][6] + A[5][6]);
  prod[1][1] <= M[1][1] * (A[1][1] + A[5][1] + A[1][5] + A[5][5]);
  prod[1][2] <= M[1][2] * (A[1][2] + A[5][2] + A[1][4] + A[5][4]);
  prod[2][0] <= M[2][0] * (A[2][0] + A[4][0] + A[2][6] + A[4][6]);
  prod[2][1] <= M[2][1] * (A[2][1] + A[4][1] + A[2][5] + A[4][5]);
  prod[2][2] <= M[2][2] * (A[2][2] + A[4][2] + A[2][4] + A[4][4]);
  prod[0][3] <= M[0][3] * (A[0][3] + A[6][3]);
  prod[1][3] <= M[1][3] * (A[1][3] + A[5][3]);
  prod[2][3] <= M[2][3] * (A[2][3] + A[4][3]);
  prod[3][0] <= M[3][0] * (A[3][0] + A[3][6]);
  prod[3][1] <= M[3][1] * (A[3][1] + A[3][5]);
  prod[3][2] <= M[3][2] * (A[3][2] + A[3][4]);
  prod[3][3] <= M[3][2] * A[3][3];
  result <= (prod[0][0] + prod[0][1] + prod[0][2] + prod[0][3]
           + prod[1][0] + prod[1][1] + prod[1][2] + prod[1][3]
           + prod[2][0] + prod[2][1] + prod[2][2] + prod[2][3]
           + prod[3][0] + prod[3][1] + prod[3][2] + prod[3][3]) >> 10;
end

/* 
always@(*) begin
 
    {M[0][0],M[0][1],M[0][2],M[0][3],M[0][4],M[0][5],M[0][6],
     M[1][0],M[1][1],M[1][2],M[1][3],M[1][4],M[1][5],M[1][6],
     M[2][0],M[2][1],M[2][2],M[2][3],M[2][4],M[2][5],M[2][6],
     M[3][0],M[3][1],M[3][2],M[3][3],M[3][4],M[3][5],M[3][6],
     M[4][0],M[4][1],M[4][2],M[4][3],M[4][4],M[4][5],M[4][6],
     M[5][0],M[5][1],M[5][2],M[5][3],M[5][4],M[5][5],M[5][6],
     M[6][0],M[6][1],M[6][2],M[6][3],M[6][4],M[6][5],M[6][6]} 
     = {32'd5, 32'd9, 32'd14, 32'd16, 32'd14, 32'd9, 32'd5,
        32'd9, 32'd18, 32'd26, 32'd29, 32'd26, 32'd18, 32'd9,
        32'd14, 32'd26, 32'd37, 32'd42, 32'd37, 32'd26, 32'd14,
        32'd16, 32'd29, 32'd42, 32'd48, 32'd42, 32'd29, 32'd16,
        32'd14, 32'd26, 32'd37, 32'd42, 32'd37, 32'd26, 32'd14,
        32'd9, 32'd18, 32'd26, 32'd29, 32'd26, 32'd18, 32'd9,
        32'd5, 32'd9, 32'd14, 32'd16, 32'd14, 32'd9, 32'd5};

    {A[0][0],A[0][1],A[0][2],A[0][3],A[0][4],A[0][5],A[0][6],
     A[1][0],A[1][1],A[1][2],A[1][3],A[1][4],A[1][5],A[1][6],
     A[2][0],A[2][1],A[2][2],A[2][3],A[2][4],A[2][5],A[2][6],
     A[3][0],A[3][1],A[3][2],A[3][3],A[3][4],A[3][5],A[3][6],
     A[4][0],A[4][1],A[4][2],A[4][3],A[4][4],A[4][5],A[4][6],
     A[5][0],A[5][1],A[5][2],A[5][3],A[5][4],A[5][5],A[5][6],
     A[6][0],A[6][1],A[6][2],A[6][3],A[6][4],A[6][5],A[6][6]} <= input_pixels;
    
    sum = 0;
    for (i=0; i<WIDTH; i++) begin
      for (j=0; j<WIDTH; j++) begin
        sum += A[i][j] * M[i][j];
       end
     end
     result = (sum >> 10);  // result = sum/(2^10) 
     
end*/

endmodule
